	// Barrier Parameters
	parameter BARR_WIDTH = 11'd76;
	parameter BARR_HEIGHT = 11'd57;
	parameter BARR0_XSTART = 11'd54;
	parameter BARR1_XSTART = BARR0_XSTART+(2*BARR_WIDTH);
	parameter BARR2_XSTART = BARR0_XSTART+(4*BARR_WIDTH);
	parameter BARR3_XSTART = BARR0_XSTART+(6*BARR_WIDTH);
	parameter BARR_BLK_SZ = 11'd19;
	parameter BARR_YSTART = 11'd340;

